`ifndef YAPP_SVH
`define YAPP_SVH

typedef uvm_config_db#(virtual yapp_if) yapp_vif_config; 
import uvm_pkg::*;
`include "yapp_packet.sv"
`include "yapp_if.sv"
`include "yapp_tx_sequencer.sv"
`include "yapp_tx_seqs.sv"
`include "yapp_tx_driver.sv"
`include "yapp_tx_monitor.sv"
`include "yapp_tx_agent.sv"
`include "yapp_env.sv"
`include "yapp_seq_lib.sv"
`include "router_virtual_sequencer.sv"
`include "router_virtual_seqs.sv"
`include "router_tb.sv"
`include "router_test_lib.sv"
`include "yapp_router.sv"
`endif //YAPP_SVH

