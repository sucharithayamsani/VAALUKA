`ifndef YAPP_SVH
`define YAPP_SVH

typedef uvm_config_db#(virtual yapp_if) yapp_vif_config; 

`include "yapp_packet.sv"
`include "yapp_tx_monitor.sv"
`include "yapp_tx_sequencer.sv"
`include "yapp_tx_seqs.sv"
`include "yapp_if.sv"
`include "yapp_tx_driver.sv"
`include "yapp_tx_agent.sv"
`include "yapp_env.sv"
`include "../tb/router_tb.sv"
`include "../tb/yapp_seq_lib.sv"
`include "../tb/router_test_lib.sv"

`endif //YAPP_SVH

